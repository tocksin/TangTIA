/*
 * PSRAM example for Sipeed Tang Nano 9K.
 * Feng Zhou, 2022
 *
 * This shows example usage of the internal PSRAM of GW1NR-9CQN88P fpga 
 * on Tang Nano 9K. It simply writes a byte 8'b10010011 to address 0, reads it 
 * back and displays the lower 6 bits on LED.
 */
library ieee;           use ieee.std_logic_1164.all;
                        use ieee.numeric_std.all;

library work;           use work.tools_pkg.all;

entity psram_top is 
    port(   sys_clk     : in sl;  --// 27 Mhz, crystal clock from board
            sys_resetn  : in sl;
            button      : in sl;   --// 0 when pressed
            led         : out slv(5 downto 0);
            oClk        : out sl;

            O_psram_ck      : out    slv(1 downto 0);
            O_psram_ck_n    : out    slv(1 downto 0);
            IO_psram_rwds   : inout  slv(1 downto 0);
            IO_psram_dq     : inout  slv(15 downto 0);
            O_psram_reset_n : out    slv(1 downto 0);
            O_psram_cs_n    : out    slv(1 downto 0)
);
end entity psram_top;

architecture rtl of psram_top is

    signal clk              : sl;           -- 74.25 Mhz master clock
    signal memory_clk       : sl;
    signal clk_d            : sl;
    signal pll_lock         : sl;

    signal wr_data          : slv(63 downto 0);
    signal rd_data          : slv(63 downto 0);
    signal rd_data_valid    : sl;
    signal addr             : slv(20 downto 0);
    signal cmd              : sl;
    signal cmd_en           : sl;
    signal data_mask        : slv(7 downto 0);

    signal state            : sl;           --// 0: write a byte, 1: read the byte back
    signal cycle            : unsigned(5 downto 0);     --// 14 cycles between write and read
    signal read_back        : slv(7 downto 0);
    signal read_count       : unsigned(7 downto 0);
    signal read_cycles      : slv(5 downto 0);
    signal testCount        : unsigned(63 downto 0);
    signal calib            : sl;
    
begin

    --// PLL to generate 148.5 Mhz memory_clk
--    Gowin_rPLL pll( .clkout(memory_clk), .lock(pll_lock), .clkoutd(clk_d), .clkin(sys_clk));
    psram_pll : entity work.Gowin_rPLL
        port map( clkin   => sys_clk,          -- 27 MHz
                  clkout  => memory_clk,       -- 50.35MHz  (50.1429)
                  clkoutd => clk_d,       -- 25.175 MHz
                  lock    => pll_lock);

-- // HS PSRAM IP (version 1, single channel)
-- // All settings are set to default, except "burst length" which is 16
-- PSRAM_Memory_Interface_HS_Top psram(
    -- .clk(sys_clk), .memory_clk(memory_clk), .pll_lock(pll_lock), .rst_n(1'b1),
    -- .O_psram_ck(O_psram_ck), .O_psram_ck_n(O_psram_ck_n), .IO_psram_rwds(IO_psram_rwds),
    -- .IO_psram_dq(IO_psram_dq), .O_psram_reset_n(O_psram_reset_n), .O_psram_cs_n(O_psram_cs_n),
    -- .addr(addr), .wr_data(wr_data), .rd_data(rd_data), .rd_data_valid(rd_data_valid),
    -- .cmd(cmd), .cmd_en(cmd_en), .data_mask(data_mask),
    -- .clk_out(clk), .init_calib(calib)
-- );
    memoryComp: entity work.PSRAM_Memory_Interface_HS_Top
        port map (
            clk             => sys_clk,             --input generated by same pll, divided by 4 normally
            memory_clk      => memory_clk,             --input usually from pll? (50-250MHz)
            --memory_clk_p    => clkFastPhased,       --input usually from pll, but phase shift 90 degrees
            pll_lock        => pll_lock,                --input use with memory clock
            rst_n           => sys_resetn,           --input active low reset

            init_calib      => calib,          --output initialization completed
            addr            => addr,           --input address (21-bit)
            wr_data         => wr_data,         --input write data (64-bit)
            data_mask       => data_mask,           --input mask for wr_data (8-bits)
            rd_data         => rd_data,         --output read data (64-bit)
            rd_data_valid   => rd_data_valid,        --output read data 1 = valid
            cmd             => cmd,             --input command channel (0=read, 1=write)
            cmd_en          => cmd_en,             --input command enable
            clk_out         => clk,              --output of 1/2 memory_clk

            -- To top level external ports
            O_psram_ck      => O_psram_ck,          -- clock
            O_psram_ck_n    => O_psram_ck_n,        -- clock inverted
            IO_psram_dq     => IO_psram_dq,         -- data in and out
            IO_psram_rwds   => IO_psram_rwds,       -- read/write control
            O_psram_cs_n    => O_psram_cs_n,        -- chip select active low
            O_psram_reset_n => O_psram_reset_n      -- reset active low
        );
  
    data_mask <= x"00";
    addr <= (others => '0');
--    wr_data <= x"00000000000000" & "01011110";
    wr_data <= slv(testCount);

    -- when button (S2 on board) is pressed, show latency in cycles
    led <= not read_back(5 downto 0) when button='1' else not read_cycles;

    process (clk, sys_resetn)
    begin
        if (sys_resetn='0') then
            state <= '0';
            cycle <= (others => '0');
            cmd_en <= '0';
            read_cycles <= (others => '0');
            read_back <= (others => '0');
        elsif rising_edge(clk) then
            -- // Read takes 22 cycles. Write takes 14
            testCount <= testCount + 1;
            cmd_en <= '0';
            
            if (calib='1') then
                cycle <= cycle + 1;
                if (state = '0') then 
                    -- write state
                    cmd <= '1';
                    if (cycle = 0) then 
                        cmd_en <= '1';  -- write enable on first cycle
                    elsif (cycle = x"C") then      -- IPUG 943 - Table 4-2, Tcmd is 14 when burst==16
                        cycle <= "000000";
                        state <= '1';          -- move to read state
                    end if;
                else
                    -- read state
                    cmd <= '0';
                    if (cycle = 0) then
                        cmd_en <= '1';  -- read enable on first cycle
                        read_count <= (others => '0');
                    else
                        if (rd_data_valid = '1') then
                            read_count <= read_count + 1;
                            if (read_count = 0) then
                                read_back <= rd_data(27 downto 20);
                            elsif (read_count = "11") then
                                read_cycles <= slv(cycle);
                                cycle <= "000000";
                                state <= '0';          -- move to write state
                            end if;
                        end if;
                    end if;
                end if;
            end if;
        end if;
    end process;

    oClk <= clk;

end architecture rtl;